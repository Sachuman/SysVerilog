
package dv_pkg;

import float_pkg::*;

import "DPI-C" function real float2real(int in);
import "DPI-C" function int real2float(real in);

function automatic float_t rand_raw_float();
    // TODO
endfunction

endpackage
