
// ## r2g





